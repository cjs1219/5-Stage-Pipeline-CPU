
module Slt(less, sum);

    input less;
    output sum;
    
    wire   sum;

    assign sum = less;

endmodule
